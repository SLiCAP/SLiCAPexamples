ModelsAndLibraries
.lib myLib.lib
.source V1
.detector V_out
.lgref E_O1
C1 out 0 C value={C_ell} vinit=0
O1 2 1 out 0 myOpAmp
R1 3 2 R value={R_s} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R2 out 1 R value={(A_v-1)*R_a} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R3 1 0 R value={R_a} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
V1 3 0 V value=0 noise=0 dc=0 dcvar=0
.end